module ila_0 (
	input logic clk,
	input logic [112:0] probe0
);

wire tmp_clk = clk;
wire [112:0] tmp_probe0 = probe0;

endmodule
